** sch_path: /home/designer/shared/OS_AnalogIC_UCLouvain_Oct2025/design_data/tb_3stage_RO.sch
**.subckt tb_3stage_RO
x1 V_2 V_1 VCC VSS sg13g2_inv_2
x2 V_3 V_2 VCC VSS sg13g2_inv_2
x3 V_1 V_3 VCC VSS sg13g2_inv_2
**** begin user architecture code

.include /opt/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
vvcc vcc 0 dc 1.2
vvss vss 0 0
.option temp = 200
.ic v(V_1) = 0
.ic v(V_2) = 1.2

.control
   tran 10p 10n
   wrdata TT_3stage_RO_v1p1.txt v(V_1)
   plot v(V_1) v(V_2) v(V_3)
.endc




.param corner=0

.if (corner==0)
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.endif

**** end user architecture code
**.ends
.end
