** sch_path: /home/designer/shared/OS_AnalogIC_VLSISOC_Oct2025/design_data/large_delay/tb_largedelay_vto1p1.sch
**.subckt tb_largedelay_vto1p1
VCC VCC GND 1.2
VSS VSS GND 0
VIN VIN VSS PULSE(0 1.2 3u 1n 1n 12u 24u)
C1 VOUT VSS 10f m=1
x1 VCC VSS VIN VOUT large_delay_vto1p1
**** begin user architecture code


.option scale=1e-6
.save v(vin) v(vout)
.control
tran 2n 6u
plot v(vin) v(vout)
plot v(vin) v(vout)+2
.endc

.measure tran tdelay
+ TRIG tran1.V(VIN) TD=0u VAL=0.6 RISE=1
+ TARG tran1.V(VOUT) TD=0u VAL=0.6 RISE=1






.param corner=0

.if (corner==0)
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
.endif

.include /opt/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**** end user architecture code
**.ends

* expanding   symbol:  large_delay_vto1p1.sym # of pins=4
** sym_path: /home/designer/shared/OS_AnalogIC_VLSISOC_Oct2025/design_data/large_delay/large_delay_vto1p1.sym
** sch_path: /home/designer/shared/OS_AnalogIC_VLSISOC_Oct2025/design_data/large_delay/large_delay_vto1p1.sch
.subckt large_delay_vto1p1 VCC VSS VIN VOUT
*.iopin VIN
*.iopin VOUT
*.iopin VCC
*.iopin VSS
x1[0] VIN VCC VSS n2 sg13g2_dlygate4sd3_1
x1[1] n2 VCC VSS n3 sg13g2_dlygate4sd3_1
x1[2] n3 VCC VSS VOUT sg13g2_dlygate4sd3_1
.ends

.GLOBAL GND
.end
